*************Decoder HSPICE netlist************ 
.include 'D:\lerning\Guilan University\VLSI\HSPICE\Low Power Full Adder - Copy\mosistsmc180.lib'
*netlist--------------------------------------- 
.global VDD GND
*-------------------------------------------------------input-------------------------------------------
VDD vdd gnd 1.8
VA0 A0 gnd 1.8
VA1 A1 gnd 1.8 
VA2 A2 gnd 1.8    
VA3 A3 gnd 1.8 
VA4 A4 gnd 1.8
VA6 Data gnd PULSE 0 1.8 .1NS 10PS 10PS 4NS 8NS
VA7 ENBB gnd 0
VA10 ENBD gnd PULSE 0 1.8 .1NS 10PS 10PS 8NS 16NS
VA8 WL gnd 0
VA9 Sen gnd PULSE 1.8 0 .1NS 10PS 10PS 16NS 32NS

*----------------------------------------------------------Inverter for decoder------------------------
.subckt Inv a ab
MIP1 vdd a ab vdd PMOS L=.18u W=.36u 
MIN1 ab a gnd gnd NMOS L=.18u W=.18u
.ends
*----------------------------------------------------------NAND2 for decoder + inv----------------------
.subckt NAND2 a b f 
MNN21 cf a 5 gnd NMOS L=.18u W=.18u
MNN22 5 b gnd gnd NMOS L=.18u W=.18u


MNP21 vdd a cf vdd PMOS L=.18u W=.36u  
MNP22 vdd b cf vdd PMOS L=.18u W=.36u

XIN cf f Inv 
.ends
*----------------------------------------------------------NAND5 for decoder + inv----------------------
.subckt NAND5 a b c d e g
XN51 a b ab NAND2
XN52 c d cd NAND2
XN53 ab cd abcd NAND2
XN54 abcd e g NAND2 
.ends
*---------------------------------------------------------SRAM Cells -----------------------------------
.subckt SRC BT BTB WL 
MSP1 vdd 3 2 vdd PMOS L=.18u W=.18u 
MSN1 2 3 gnd gnd NMOS L=.18u W=.62u

MSP2 vdd 2 3 vdd PMOS L=.18u W=.28u  
MSN2 3 2 gnd gnd NMOS L=.18u W=.82u

MSN3 BT WL 2 gnd NMOS L=.18u W=.36u
MSN4 BTB WL 3 gnd NMOS L=.18u W=.36u

C1 BT 0 10f
C2 BTB 0 10f
.ends
*-------------------------------------------------------BTline Conditional--------------------------------------------------------------------------
.subckt BTCL ENBB BTN BTBN
MBTP1 vdd ENBB BTN vdd PMOS L=.18u W=.63u
MBTP2 vdd ENBB BTBN vdd PMOS L=.18u W=.63u
.ends
*-------------------------------------------------------Read Circuit-------------------------------------------------------------------
.subckt RDC ENBB BTN BTBN OUTBTN OUTBTBN
*XBTLRDC ENBB BTN BTBN BTCL
XIRC1 BTN OUTBTN Inv
XIRC2 BTBN OUTBTBN Inv
.ends
*-------------------------------------------------------WRITE Circuit-------------------------------------------------------------------------
.subckt WRC ENBB WL Data BTN BTBN
XI1 data datab Inv

MWRN1 BTN WL W1 gnd NMOS L=.18u W=.82u
MWRN2 W1 Datab gnd gnd NMOS L=.18u W=.82u

MWRN3 BTBN WL W2 gnd NMOS L=.18u W=.82u
MWRN4 W2 Data gnd gnd NMOS L=.18u W=.82u
.ends
*-------------------------------------------------------Sense--------------------------------------------------------------
*.subckt Sense BTN BTBN Sen DataS DatabS 
*XSI3 Sen Senb Inv

*MSEP6 BTBN Senb 24 vdd PMOS L=.18u W=.72u 

*MSEP24 vdd 13 24 vdd PMOS L=.18u W=.72u 
*MSEN24 24 13 1324 gnd NMOS L=.18u W=.36u


*MSEP13 vdd 24 13 vdd PMOS L=.18u W=.72u  
*MSEN13 13 24 1324 gnd NMOS L=.18u W=.36u

*MSEP5 BTN Senb 13 vdd PMOS L=.18u W=.72u

*MSEN7 1324 24 gnd gnd NMOS L=.18u W=.36u

*XSI1 24 databS Inv
*XSI2 13 dataS Inv

*.ends
*---------------------------------------------------------Decoder5*32-----------------------------------
.subckt DCR5 A0 A1 A2 A3 A4 ENBD D0 D1 D2 D3 D4 D5 D6 D7 D8 D9 D10 D11 D12 D13 D14 D15 D16 D17 D18 D19 D20 D21 D22 D23 D24 D25 D26 D27 D28 D29 D30 D31
XI0 A0 A0B Inv
XI1 A1 A1B Inv
XI2 A2 A2B Inv
XI3 A3 A3B Inv
XI4 A4 A4B Inv

XNDCR0 A0B A1B A2B A3B A4B Dn0 NAND5
XNDCR1 A0B A1B A2B A3B A4 Dn1 NAND5
XNDCR2 A0B A1B A2B A3 A4B Dn2 NAND5
XNDCR3 A0B A1B A2B A3 A4 Dn3 NAND5
XNDCR4 A0B A1B A2 A3B A4B Dn4 NAND5
XNDCR5 A0B A1B A2 A3B A4 Dn5 NAND5
XNDCR6 A0B A1B A2 A3 A4B Dn6 NAND5
XNDCR7 A0B A1B A2 A3 A4 Dn7 NAND5
XNDCR8 A0B A1 A2B A3B A4B Dn8 NAND5
XNDCR9 A0B A1 A2B A3B A4 Dn9 NAND5
XNDCR10 A0B A1 A2B A3 A4B Dn10 NAND5
XNDCR11 A0B A1 A2B A3 A4 Dn11 NAND5
XNDCR12 A0B A1 A2 A3B A4B Dn12 NAND5
XNDCR13 A0B A1 A2 A3B A4 Dn13 NAND5
XNDCR14 A0B A1 A2 A3 A4B Dn14 NAND5
XNDCR15 A0B A1 A2 A3 A4 Dn15 NAND5
XNDCR16 A0 A1B A2B A3B A4B Dn16 NAND5
XNDCR17 A0 A1B A2B A3B A4 Dn17 NAND5
XNDCR18 A0 A1B A2B A3 A4B Dn18 NAND5
XNDCR19 A0 A1B A2B A3 A4 Dn19 NAND5
XNDCR20 A0 A1B A2 A3B A4B Dn20 NAND5
XNDCR21 A0 A1B A2 A3B A4 Dn21 NAND5
XNDCR22 A0 A1B A2 A3 A4B Dn22 NAND5
XNDCR23 A0 A1B A2 A3 A4 Dn23 NAND5
XNDCR24 A0 A1 A2B A3B A4B Dn24 NAND5
XNDCR25 A0 A1 A2B A3B A4 Dn25 NAND5
XNDCR26 A0 A1 A2B A3 A4B Dn26 NAND5
XNDCR27 A0 A1 A2B A3 A4 Dn27 NAND5
XNDCR28 A0 A1 A2 A3B A4B Dn28 NAND5
XNDCR29 A0 A1 A2 A3B A4 Dn29 NAND5
XNDCR30 A0 A1 A2 A3 A4B Dn30 NAND5
XNDCR31 A0 A1 A2 A3 A4 Dn31 NAND5

XN20 Dn0 ENBD D0 NAND2
XN21 Dn1 ENBD D1 NAND2
XN22 Dn2 ENBD D2 NAND2
XN23 Dn3 ENBD D3 NAND2
XN24 Dn4 ENBD D4 NAND2
XN25 Dn5 ENBD D5 NAND2
XN26 Dn6 ENBD D6 NAND2
XN27 Dn7 ENBD D7 NAND2
XN28 Dn8 ENBD D8 NAND2
XN29 Dn9 ENBD D9 NAND2
XN210 Dn10 ENBD D10 NAND2
XN211 Dn11 ENBD D11 NAND2
XN212 Dn12 ENBD D12 NAND2
XN213 Dn13 ENBD D13 NAND2
XN214 Dn14 ENBD D14 NAND2
XN215 Dn15 ENBD D15 NAND2
XN216 Dn16 ENBD D16 NAND2
XN217 Dn17 ENBD D17 NAND2
XN218 Dn18 ENBD D18 NAND2
XN219 Dn19 ENBD D19 NAND2
XN220 Dn20 ENBD D20 NAND2
XN221 Dn21 ENBD D21 NAND2
XN222 Dn22 ENBD D22 NAND2
XN223 Dn23 ENBD D23 NAND2
XN224 Dn24 ENBD D24 NAND2
XN225 Dn25 ENBD D25 NAND2
XN226 Dn26 ENBD D26 NAND2
XN227 Dn27 ENBD D27 NAND2
XN228 Dn28 ENBD D28 NAND2
XN229 Dn29 ENBD D29 NAND2
XN230 Dn30 ENBD D30 NAND2
XN231 Dn31 ENBD D31 NAND2
.ends

*-------------------------------------------------------SRAM Column UNIT------------------------------------------------------------------------
.subckt SRU BTN0 BTN1 BTN2 BTN3 BTN4 BTN5 BTN6 BTN7 BTN8 BTN9 BTN10 BTN11 BTN12 BTN13 BTN14 BTN15 BTN16 BTN17 BTN18 BTN19 BTN20 BTN21 BTN22 BTN23 BTN24 BTN25 BTN26 BTN27 BTN28 BTN29 BTN30 BTN31 BTBN0 BTBN1 BTBN2 BTBN3 BTBN4 BTBN5 BTBN6 BTBN7 BTBN8 BTBN9 BTBN10 BTBN11 BTBN12 BTBN13 BTBN14 BTBN15 BTBN16 BTBN17 BTBN18 BTBN19 BTBN20 BTBN21 BTBN22 BTBN23 BTBN24 BTBN25 BTBN26 BTBN27 BTBN28 BTBN29 BTBN30 BTBN31 D0 D1 D2 D3 D4 D5 D6 D7 D8 D9 D10 D11 D12 D13 D14 D15 D16 D17 D18 D19 D20 D21 D22 D23 D24 D25 D26 D27 D28 D29 D30 D31 Data WL OUTBTN OUTBTBN

XSRU1 BTN0 BTBN0 D0 SRC
R1 BTN0 BTN1 10
R2 BTBN0 BTBN1 10 
XSRU2 BTN1 BTBN D1 SRC
R3 BTN1 BTN2 10
R4 BTBN1 BTBN2 10 
XSRU3 BTN2 BTBN2 D2 SRC
R5 BTN2 BTN3 10
R6 BTBN2 BTBN3 10 
XSRU4 BTN3 BTBN3 D3 SRC
R7 BTN3 BTN4 10
R8 BTBN3 BTBN4 10 
XSRU5 BTN4 BTBN4 D4 SRC
R9 BTN4 BTN5 10
R10 BTBN4 BTBN5 10
XSRU6 BTN5 BTBN5 D5 SRC
R11 BTN5 BTN6 10
R12 BTBN5 BTBN6 10
XSRU7 BTN6 BTBN6 D6 SRC
R13 BTN6 BTN7 10
R14 BTBN6 BTBN7 10
XSRU8 BTN7 BTBN7 D7 SRC
R15 BTN7 BTN8 10
R16 BTBN7 BTBN8 10
XSRU9 BTN8 BTBN8 D8 SRC
R17 BTN8 BTN9 10
R18 BTBN8 BTBN9 10
XSRU10 BTN9 BTBN9 D9 SRC
R19 BTN9 BTN10 10
R20 BTBN9 BTBN10 10
XSRU11 BTN10 BTBN10 D10 SRC
R21 BTN10 BTN11 10
R22 BTBN10 BTBN11 10
XSRU12 BTN11 BTBN11 D11 SRC
R23 BTN11 BTN12 10
R24 BTBN11 BTBN12 10
XSRU13 BTN12 BTBN12 D12 SRC
R25 BTN12 BTN13 10
R26 BTBN12 BTBN13 10
XSRU14 BTN13 BTBN13 D13 SRC
R27 BTN13 BTN14 10
R28 BTBN13 BTBN14 10
XSRU15 BTN14 BTBN14 D14 SRC
R29 BTN14 BTN15 10
R30 BTBN14 BTBN15 10
XSRU16 BTN15 BTBN15 D15 SRC
R31 BTN15 BTN16 10
R32 BTBN15 BTBN16 10
XSRU17 BTN16 BTBN16 D16 SRC
R33 BTN16 BTN17 10
R34 BTBN16 BTBN17 10
XSRU18 BTN17 BTBN17 D17 SRC
R35 BTN17 BTN18 10
R36 BTBN17 BTBN18 10
XSRU19 BTN18 BTBN18 D18 SRC
R37 BTN18 BTN19 10
R38 BTBN18 BTBN19 10
XSRU20 BTN19 BTBN19 D19 SRC
R39 BTN19 BTN20 10
R40 BTBN19 BTBN20 10
XSRU21 BTN20 BTBN20 D20 SRC
R41 BTN20 BTN21 10
R42 BTBN20 BTBN21 10
XSRU22 BTN21 BTBN21 D21 SRC
R43 BTN21 BTN22 10
R44 BTBN21 BTBN22 10
XSRU23 BTN22 BTBN22 D22 SRC
R45 BTN22 BTN23 10
R46 BTBN22 BTBN23 10
XSRU24 BTN23 BTBN23 D23 SRC
R47 BTN23 BTN24 10
R48 BTBN23 BTBN24 10
XSRU25 BTN24 BTBN24 D24 SRC
R49 BTN24 BTN25 10
R50 BTBN24 BTBN25 10
XSRU26 BTN25 BTBN25 D25 SRC
R51 BTN25 BTN26 10
R52 BTBN25 BTBN26 10
XSRU27 BTN26 BTBN26 D26 SRC
R53 BTN26 BTN27 10
R54 BTBN26 BTBN27 10
XSRU28 BTN27 BTBN27 D27 SRC
R55 BTN27 BTN28 10
R56 BTBN27 BTBN28 10
XSRU29 BTN28 BTBN28 D28 SRC
R57 BTN28 BTN29 10
R58 BTBN28 BTBN29 10
XSRU30 BTN29 BTBN29 D29 SRC
R59 BTN29 BTN30 10
R60 BTBN29 BTBN30 10
XSRU31 BTN30 BTBN30 D30 SRC
R61 BTN30 BTN31 10
R62 BTBN30 BTBN31 10
XSRU32 BTN31 BTBN31 D31 SRC

XBTLRDC ENBB BTN0 BTBN0 BTCL
*XSEN1 BTN31 BTBN31 Sen DataS DatabS Sense
XRDC1 ENBB BTN31 BTBN31 OUTBTN OUTBTBN RDC
XWRC1 ENBB WL Data BTN31 BTBN31 WRC

.ends
*-------------------------------------------------------SRAM 32*8------------------------------------------------------------------------------
XDC1 A0 A1 A2 A3 A4 ENBD D0 D1 D2 D3 D4 D5 D6 D7 D8 D9 D10 D11 D12 D13 D14 D15 D16 D17 D18 D19 D20 D21 D22 D23 D24 D25 D26 D27 D28 D29 D30 D31 DCR5

XSRR0 BT0 BT01 BT02 BT03 BT04 BT05 BT06 BT07 BT08 BT09 BT010 BT011 BT012 BT013 BT014 BT015 BT016 BT017 BT018 BT019 BT020 BT021 BT022 BT023 BT024 BT025 BT026 BT027 BT028 BT029 BT030 BT031 BTB0 BTB01 BTB02 BTB03 BTB04 BTB05 BTB06 BTB07 BTB08 BTB09 BTB010 BTB011 BTB012 BTB013 BTB014 BTB015 BTB016 BTB017 BTB018 BTB019 BTB020 BTB021 BTB022 BTB023 BTB024 BTB025 BTB026 BTB027 BTB028 BTB029 BTB030 BTB031 D0 D1 D2 D3 D4 D5 D6 D7 D8 D9 D10 D11 D12 D13 D14 D15 D16 D17 D18 D19 D20 D21 D22 D23 D24 D25 D26 D27 D28 D29 D30 D31 Data WL OUTBT0 OUTBTB0 SRU
XSRR1 BT1 BT11 BT12 BT13 BT14 BT15 BT16 BT17 BT18 BT19 BT110 BT111 BT112 BT113 BT114 BT115 BT116 BT117 BT118 BT119 BT120 BT121 BT122 BT123 BT124 BT125 BT126 BT127 BT128 BT129 BT130 BT131 BTB1 BTB11 BTB12 BTB13 BTB14 BTB15 BTB16 BTB17 BTB18 BTB19 BTB110 BTB111 BTB112 BTB113 BTB114 BTB115 BTB116 BTB117 BTB118 BTB119 BTB120 BTB121 BTB122 BTB123 BTB124 BTB125 BTB126 BTB127 BTB128 BTB129 BTB130 BTB131 D0 D1 D2 D3 D4 D5 D6 D7 D8 D9 D10 D11 D12 D13 D14 D15 D16 D17 D18 D19 D20 D21 D22 D23 D24 D25 D26 D27 D28 D29 D30 D31 Data WL OUTBT1 OUTBTB1 SRU
XSRR2 BT2 BT21 BT22 BT23 BT24 BT25 BT26 BT27 BT28 BT29 BT210 BT211 BT212 BT213 BT214 BT215 BT216 BT217 BT218 BT219 BT220 BT221 BT222 BT223 BT224 BT225 BT226 BT227 BT228 BT229 BT230 BT231 BTB2 BTB21 BTB22 BTB23 BTB24 BTB25 BTB26 BTB27 BTB28 BTB29 BTB210 BTB211 BTB212 BTB213 BTB214 BTB215 BTB216 BTB217 BTB218 BTB219 BTB220 BTB221 BTB222 BTB223 BTB224 BTB225 BTB226 BTB227 BTB228 BTB229 BTB230 BTB231 D0 D1 D2 D3 D4 D5 D6 D7 D8 D9 D10 D11 D12 D13 D14 D15 D16 D17 D18 D19 D20 D21 D22 D23 D24 D25 D26 D27 D28 D29 D30 D31 Data WL OUTBT2 OUTBTB2 SRU
XSRR3 BT3 BT31 BT32 BT33 BT34 BT35 BT36 BT37 BT38 BT39 BT310 BT311 BT312 BT313 BT314 BT315 BT316 BT317 BT318 BT319 BT320 BT321 BT322 BT323 BT324 BT325 BT326 BT327 BT328 BT329 BT330 BT331 BTB3 BTB31 BTB32 BTB33 BTB34 BTB35 BTB36 BTB37 BTB38 BTB39 BTB310 BTB311 BTB312 BTB313 BTB314 BTB315 BTB316 BTB317 BTB318 BTB319 BTB320 BTB321 BTB322 BTB323 BTB324 BTB325 BTB326 BTB327 BTB328 BTB329 BTB330 BTB331 D0 D1 D2 D3 D4 D5 D6 D7 D8 D9 D10 D11 D12 D13 D14 D15 D16 D17 D18 D19 D20 D21 D22 D23 D24 D25 D26 D27 D28 D29 D30 D31 Data WL OUTBT3 OUTBTB3 SRU
XSRR4 BT4 BT41 BT42 BT43 BT44 BT45 BT46 BT47 BT48 BT49 BT410 BT411 BT412 BT413 BT414 BT415 BT416 BT417 BT418 BT419 BT420 BT421 BT422 BT423 BT424 BT425 BT426 BT427 BT428 BT429 BT430 BT431 BTB4 BTB41 BTB42 BTB43 BTB44 BTB45 BTB46 BTB47 BTB48 BTB49 BTB410 BTB411 BTB412 BTB413 BTB414 BTB415 BTB416 BTB417 BTB418 BTB419 BTB420 BTB421 BTB422 BTB423 BTB424 BTB425 BTB426 BTB427 BTB428 BTB429 BTB430 BTB431 D0 D1 D2 D3 D4 D5 D6 D7 D8 D9 D10 D11 D12 D13 D14 D15 D16 D17 D18 D19 D20 D21 D22 D23 D24 D25 D26 D27 D28 D29 D30 D31 Data WL OUTBT4 OUTBTB4 SRU
XSRR5 BT5 BT51 BT52 BT53 BT54 BT55 BT56 BT57 BT58 BT59 BT510 BT511 BT512 BT513 BT514 BT515 BT516 BT517 BT518 BT519 BT520 BT521 BT522 BT523 BT524 BT525 BT526 BT527 BT528 BT529 BT530 BT531 BTB5 BTB51 BTB52 BTB53 BTB54 BTB55 BTB56 BTB57 BTB58 BTB59 BTB510 BTB511 BTB512 BTB513 BTB514 BTB515 BTB516 BTB517 BTB518 BTB519 BTB520 BTB521 BTB522 BTB523 BTB524 BTB525 BTB526 BTB527 BTB528 BTB529 BTB530 BTB531 D0 D1 D2 D3 D4 D5 D6 D7 D8 D9 D10 D11 D12 D13 D14 D15 D16 D17 D18 D19 D20 D21 D22 D23 D24 D25 D26 D27 D28 D29 D30 D31 Data WL OUTBT5 OUTBTB5 SRU 
XSRR6 BT6 BT61 BT62 BT63 BT64 BT65 BT66 BT67 BT68 BT69 BT610 BT611 BT612 BT613 BT614 BT615 BT616 BT617 BT618 BT619 BT620 BT621 BT622 BT623 BT624 BT625 BT626 BT627 BT628 BT629 BT630 BT631 BTB6 BTB61 BTB62 BTB63 BTB64 BTB65 BTB66 BTB67 BTB68 BTB69 BTB610 BTB611 BTB612 BTB613 BTB614 BTB615 BTB616 BTB617 BTB618 BTB619 BTB620 BTB621 BTB622 BTB623 BTB624 BTB625 BTB626 BTB627 BTB628 BTB629 BTB630 BTB631 D0 D1 D2 D3 D4 D5 D6 D7 D8 D9 D10 D11 D12 D13 D14 D15 D16 D17 D18 D19 D20 D21 D22 D23 D24 D25 D26 D27 D28 D29 D30 D31 Data WL OUTBT6 OUTBTB6 SRU
XSRR7 BT7 BT71 BT72 BT73 BT74 BT75 BT76 BT77 BT78 BT79 BT710 BT711 BT712 BT713 BT714 BT715 BT716 BT717 BT718 BT719 BT720 BT721 BT722 BT723 BT724 BT725 BT726 BT727 BT728 BT729 BT730 BT731 BTB7 BTB71 BTB72 BTB73 BTB74 BTB75 BTB76 BTB77 BTB78 BTB79 BTB710 BTB711 BTB712 BTB713 BTB714 BTB715 BTB716 BTB717 BTB718 BTB719 BTB720 BTB721 BTB722 BTB723 BTB724 BTB725 BTB726 BTB727 BTB728 BTB729 BTB730 BTB731 D0 D1 D2 D3 D4 D5 D6 D7 D8 D9 D10 D11 D12 D13 D14 D15 D16 D17 D18 D19 D20 D21 D22 D23 D24 D25 D26 D27 D28 D29 D30 D31 Data WL OUTBT7 OUTBTB7 SRU


*-------------------------------------------------------TRAN-------------------------------------------------------------------------------------

.options post=2 nomod 
.op 
.TRAN 1ps 32ns * transient analysis: Step end_time 
.end